Computation test

ADDI X10, XZR, 10

1001 0001 0000 0000 0010 1000 0000 01010

ADDI X11, XZR, 8

1001 0001 0000 0000 0010 0000 0000 01011

ADDI X9, XZR, 100

1001 0001 0000 0001 1001 0000 0000 01001

SUBI X9, X9, 10

1101 0001 0000 0000 0010 1001 0010 1001

ADD  X10, X9, X11

1000 1011 0000 1011 0000 0001 0010 1010


Communication test

LDUR X10, [X11, 0]

1111 1000 0100 0000 0000 0001 0110 1010

STUR X10, [X9, 0]

1111 1000 0000 0000 0000 0001 0010 1010


Final test

ADDI X9, XZR, 100

1001 0001 0000 0001 1001 0000 0000 01001

SUBI X9, X9, 1

1101 0001 0000 0000 0000 0101 0010 1001

ADDI X11, X11, 8

1001 0001 0000 0000 0010 0001 0110 1011

ADD  X10,X9,X11

1000 1011 0000 1011 0000 0001 0010 1010

LDUR X10, [X11, 0]

11111000010 000000000 00 01011 01010

STUR X10, [X9, 0]

11111000000 000000000 00 01001 01010

CBZ X9, 4

1011 0100 0000000000000000100 01001


B l1 --7

100101 00000000000000000000000111


















